module top;
  initial begin
    run_test("test");
  end
endmodule
